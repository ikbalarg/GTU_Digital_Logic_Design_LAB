module tb_problem2();
	logic Cin,A0,B0,A1,B1,A2,B2,A3,B3,A4,B4;
	logic S0,S1,S2,S3,S4,Cout;
problem2 dut0(Cin,A0,B0,A1,B1,A2,B2,A3,B3,A4,B4,S0,S1,S2,S3,S4,Cout);
initial begin
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=0;A3=0;B3=0;A4=0;B4=0;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=0;A3=0;B3=0;A4=0;B4=1;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=0;A3=0;B3=0;A4=1;B4=1;#10
	Cin=1;A0=0;B0=1;A1=0;B1=1;A2=0;B2=0;A3=0;B3=0;A4=1;B4=0;#10
	Cin=0;A0=1;B0=1;A1=0;B1=0;A2=0;B2=0;A3=0;B3=0;A4=0;B4=0;#10
	Cin=1;A1=0;B0=1;A1=0;B1=0;A2=0;B2=0;A3=0;B3=0;A4=0;B4=0;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=0;A3=0;B3=1;A4=1;B4=1;#10
	Cin=0;A0=0;B0=1;A1=0;B1=0;A2=0;B2=0;A3=1;B3=1;A4=1;B4=1;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=1;A3=1;B3=0;A4=0;B4=0;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=1;A3=1;B3=1;A4=1;B4=0;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=0;B2=1;A3=1;B3=1;A4=1;B4=1;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=1;B2=1;A3=0;B3=0;A4=0;B4=0;#10
	Cin=0;A0=0;B0=0;A1=0;B1=0;A2=1;B2=1;A3=0;B3=1;A4=1;B4=0;#10
	Cin=1;A0=0;B0=0;A1=0;B1=1;A2=0;B2=0;A3=0;B3=0;A4=0;B4=0;#10
	Cin=1;A0=0;B0=0;A1=0;B1=0;A2=0;B2=0;A3=1;B3=1;A4=1;B4=1;#10
	Cin=1;A0=1;B0=1;A1=1;B1=1;A2=1;B2=1;A3=1;B3=1;A4=1;B4=1;#10
	$stop;
  end
endmodule
